`define ALU_ADD 3'b000
`define ALU_SUB 3'b001
`define ALU_AND 3'b010
`define ALU_OR  3'b011
`define ALU_XOR 3'b100
`define ALU_SLT 3'b101
`define ALU_SL  3'b110
`define ALU_SR  3'b111
`define ALU_DCR 3'bxxx
